** Profile: "SCHEMATIC1-test"  [ C:\Users\29721\Desktop\prectice\test-pspicefiles\schematic1\test.sim ] 

** Creating circuit file "test.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "C:/Cadence/Cadence_SPB_16.6-2015/tools/pspice/library/STGW40H65DFB-V2.lib" 
* From [PSPICE NETLIST] section of C:\Cadence\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 
.lib "C:\Cadence\Cadence_SPB_16.6-2015\tools\capture\library\pspice\STGW40H65DFB-V2.OLB" 

*Analysis directives: 
.TRAN  0 0.08 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
